//-----------------------------------------------------
// Design Name : ram_dp_ar_aw
// File Name   : ram_dp_ar_aw.v
// Function    : Asynchronous read write RAM
// Coder       : Deepak Kumar Tala
//-----------------------------------------------------
module ram_dp_ar_aw(
address_0 , // address_0 Input
data_0    , // data_0 bi-directional
cs_0      , // Chip Select
we_0      , // Write Enable/Read Enable
address_1 , // address_1 Input
data_1    , // data_1 bi-directional
cs_1      , // Chip Select
we_1      , // Write Enable/Read Enable
oe_1        // Output Enable
); 

	parameter DATA_WIDTH = 12;
	parameter ADDR_WIDTH = 3 ;
	parameter RAM_DEPTH = 8;

	//--------------Input Ports----------------------- 
	input [ADDR_WIDTH-1:0] address_0 ;
	input cs_0 ;
	input we_0 ;
	input [ADDR_WIDTH-1:0] address_1 ;
	input cs_1 ;
	input we_1 ;
	input oe_1 ; 

	//--------------Inout Ports----------------------- 
	input [DATA_WIDTH-1:0] data_0 ; 
	output [DATA_WIDTH-1:0] data_1 ;

	//--------------Internal variables---------------- 
	//reg [DATA_WIDTH-1:0] data_0_out ; 
	reg [DATA_WIDTH-1:0] data_1_out ;
	reg [DATA_WIDTH-1:0] mem [0:RAM_DEPTH-1];


	//--------------Code Starts Here------------------ 
	// Memory Write Block 
	// Write Operation : When we_0 = 1, cs_0 = 1

	always @ (address_0 or cs_0 or we_0 or data_0)
	begin : MEM_WRITE
		if ( cs_0 && we_0 ) begin
			 mem[address_0] = data_0;
		end
		//else if  (cs_1 && we_1) begin
		//	 mem[address_1] = data_1;
		//end
	end

	assign data_1 = data_1_out;
	// Memory Read Block 1 
	// Read Operation : When we_1 = 0, oe_1 = 1, cs_1 = 1
	always @ (address_1 or cs_1 or we_1 or oe_1)
	begin : MEM_READ_1
		if (cs_1 && !we_1 && oe_1) begin
			data_1_out = mem[address_1]; 
		end else begin
			data_1_out = 0; 
		end
	end

endmodule // End of Module ram_dp_ar_aw

